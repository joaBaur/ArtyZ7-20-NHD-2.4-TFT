-- Company: Baur 3.0 Service GmbH
-- Engineer: Joachim Baur
-- 
-- Create Date: 01.06.2018
-- Module Name: VideoProcessing - Behavioral
-- Description: Writes video pixel data to block ram
-- video rgb data is received from dvi2rgb ip
----------------------------------------------------------------------------------

library IEEE;
use IEEE.STD_LOGIC_1164.ALL;
use IEEE.STD_LOGIC_ARITH.ALL; -- used for calculating bram_addra

entity VideoProcessing is
	Port (
		i_pxl_clock	 : in STD_LOGIC;						-- pixel clock generated by HDMI decoder
		i_rgb 		 : in STD_LOGIC_VECTOR (23 downto 0); 	-- rgb data (ordered r-b-g!)
		i_h_sync 	 : in STD_LOGIC;						-- horizontal sync signal
		i_v_sync 	 : in STD_LOGIC;						-- vertical sync signal
		i_vde 		 : in STD_LOGIC;						-- pixel data active signal

		i_resolution : in STD_LOGIC;						-- state of hardware switch SW0 
		
		bram_addra 	 : out std_logic_vector (16 downto 0);	-- adress lines of block ram port a
		bram_dina 	 : out std_logic_vector (23 downto 0);  -- data lines of block ram port a
		bram_wea 	 : out std_logic						-- write enable line of block ram port a
	);
end VideoProcessing;

architecture Behavioral of VideoProcessing is

-- registers for storing the values from the previous clock cycle
signal last_vsync : STD_LOGIC := '0';
signal last_vde   : STD_LOGIC := '0';

begin

	video_processing: process(i_pxl_clock)
	
	-- horizontal start of the 320x240 area to grab
	-- max value = 1920 - 320 = 1600 (for 1920 x 1080 resolution)
	constant h_start  : integer range 0 to 1600 := 0; 
	
	-- vertical start of the 320x240 area to grab
    -- max value = 1080 - 240 = 840 (for 1920 x 1080 resolution)
	constant v_start  : integer range 0 to  840 := 0;

	variable h_count  : integer range 0 to 1920 := 0;
    variable v_count  : integer range 0 to 1080 := 0;
    variable curr_col : integer range 0 to 1920 := 0;
    variable curr_row : integer range 0 to 1080 := 0;
    
    variable startNewFrame : STD_LOGIC := '1'; -- flag for the start of a new frame
    variable ram_address : integer range 0 to 76800 := 0;
    
	begin
		if rising_edge(i_pxl_clock) then
		
		    -- i_vde = '1': i_rgb contains pixel data (r-b-g)
		    -- i_vde = '0': i_rgb contains other/non-pixel data (blanking)

		    -- i_vde 1->0: end of a row of pixel data reached, start blanking
	        if i_vde = '0' and last_vde = '1' then
	           -- increment the row number
	           v_count := v_count + 1;
	        end if;
		   
		    -- i_v_sync 0->1: start of new frame   
		    if i_v_sync = '1' and last_vsync = '0' then
		    	-- just set the flag for the start of a new frame
		    	-- wait for i_vde to become '1' for resetting v_count
		        startNewFrame := '1';
		    end if;
		   
		    -- i_vde 0->1: new pixels start arriving (new row and maybe new frame)
		    if i_vde = '1' then
		        if last_vde = '0' then
		    	    -- reset column number to 0
		            h_count := 0;
		            if startNewFrame = '1' then
                        -- start new frame, clear flag and reset row number to 0
                        startNewFrame := '0';
                        v_count := 0;
                    end if;
		        else
		    	    -- i_de is 1, so pixel data is still arriving, increase column number
		            h_count := h_count + 1;
		        end if;
		    end if;

		    -- save values for comparison in next clock cycle
		    last_vsync <= i_v_sync;
		    last_vde   <= i_vde;
		   
		   	-- scale resolution by half if switch "i_resolution" is ON
            if i_resolution = '1' then
                curr_col := h_count/2;
                curr_row := v_count/2;
            else
                curr_col := h_count;
                curr_row := v_count;
            end if;

		    -- if the pixel data is within the tft bounds, store it in block ram
		    if curr_col >= h_start and curr_col < (h_start+320) and curr_row >= v_start and curr_row < (v_start + 240) then
		    
	            -- calculate the block ram index address
	            ram_address := (curr_row - v_start) * 320 + (curr_col - h_start);    
	                   
	            bram_addra <= conv_std_logic_vector(ram_address, bram_addra'length);
                bram_dina <= i_rgb;
                bram_wea <= '1';
	     	else 
	     		bram_wea <= '0'; -- no ram write
			end if; 
   
		end if;
	end process video_processing;

end Behavioral;